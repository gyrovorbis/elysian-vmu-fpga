
use work.memBus.all;

entity VmuLcdc is 
	port (
		memBusIn	: in VmuMemoryBusIn;
		memBusOut	: out VmuMemoryBusOut
	);

end entity;

architecture rtl of VmuLcdc is
begin

end architecture;