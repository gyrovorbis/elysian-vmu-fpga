
use work.memBus.all;

entity VmuFlash is 
	port (
		memBusIn	: in VmuMemoryBusIn;
		memBusOut	: out VmuMemoryBusOut
	);

end entity;


architecture rtl of VmuFlash is 
begin

end architecture;