
use work.memBus.all;

entity VmuRom is 
	port (
		memBusIn	: in VmuMemoryBusIn;
		memBusOut	: out VmuMemoryBusOut
	);

end entity;

architecture rtl of VMURom is 
begin

end architecture;